library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 

entity fsm_counter is 
    port(); 
end entity; 

architecture bhv of fsm_counter is 
    begin 









    end bhv; 